.title KiCad schematic
Q1 Net-_Q1-Pad1_ Net-_Q1-Pad2_ Net-_Q1-Pad3_ BC108
U1 Net-_Q1-Pad2_ Net-_Q1-Pad3_ Net-_R1-Pad1_ 7400
R1 Net-_R1-Pad1_ Net-_Q1-Pad1_ R
.end

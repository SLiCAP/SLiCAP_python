EKV model
.lib CMOS18.lib
X1 D G S 0 CMOS18P W={W} L={L} ID={-I_D} 
.param I_D=0 W=2.2e-07 L=1.8e-07
.end

ACcoupling
.detector V_out
C1 2 out C value={C_c} vinit=0
R1 2 1 R value={R_s} noisetemp=0 noiseflow=0 dcvar=0 dcvarlot=0
R2 B out R value={R_a} noisetemp=0 noiseflow=0 dcvar=0 dcvarlot=0
R3 out 0 R value={R_b} noisetemp=0 noiseflow=0 dcvar=0 dcvarlot=0
V1 B 0 V value={V_B/s} noise=0 dc=0 dcvar=0
V2 1 0 V value={V_p*2*pi*f_s/(s^2+(2*pi*f_s)^2)} noise=0 dc=0 dcvar=0
.end
"myPassiveNetwork"
.param R_a=10 G_0=1m R_b=100 R_c=2k R_d=50 L=1m C_a=1u R_b=100 C_b=1n tau=10u
.detector V_1 V_2
.source V1
C1 4 1 C value={C_a} vinit=0
C2 2 0 C value={C_b} vinit=0
G1 3 0 6 5 G value={G_0/(1+s*tau)}
L1 6 1 L value={L} iinit=0
R1 6 5 R value={R_a} noisetemp={T} noiseflow=0 dcvar={sigma_R1^2} dcvarlot=0
R2 0 2 R value={R_b} noisetemp={T} noiseflow=0 dcvar={sigma_R1^2} dcvarlot=0
R3 0 3 R value={R_c} noisetemp={T} noiseflow=0 dcvar={sigma_R1^2} dcvarlot=0
R4 0 4 R value={R_d} noisetemp={T} noiseflow=0 dcvar={sigma_R1^2} dcvarlot=0
V1 5 0 V value=0 noise={S_v} dc={V_DC} dcvar={(sigma_V*V_DC)^2}
.end
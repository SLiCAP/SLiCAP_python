"Balanced Noisy Network"
.detector V_outP V_outN
C1 outN outP C value={C_a} vinit=0
C2 0 1 C value={C_b} vinit=0
E1 CM 3 outP 0 E value=0.5
E2 3 0 outN 0 E value=0.5
I1 0 1 I value={I_s} noise={S_i} dc=0 dcvar=0
R1N inN outN R value={R_a} noisetemp={T} noiseflow=0 dcvar=0 dcvarlot=0
R1P inP outP R value={R_a} noisetemp={T} noiseflow=0 dcvar=0 dcvarlot=0
R2N outN 2 R value={R_b} noisetemp={T} noiseflow=0 dcvar=0 dcvarlot=0
R2P outP 2 R value={R_b} noisetemp={T} noiseflow=0 dcvar=0 dcvarlot=0
R3 2 0 R value={R_c} noisetemp={T} noiseflow=0 dcvar=0 dcvarlot=0
V1N inN 1 V value={V_b} noise={S_vb} dc=0 dcvar=0
V1P inP 1 V value={V_a} noise={S_va} dc=0 dcvar=0
.end
"Balanced Vamp"
.param R_a=100k R_b=100 R_s=1k R_L=200
.source V1P V1N
.detector V_outP V_outN
.param Lot_1={sigma_L^2}
E1 comm 1 outP 0 E value=0.5
E2 1 0 outN 0 E value=0.5
R1N inN srcN R value={R_s} noisetemp=0 noiseflow=0 dcvar=0 dcvarlot=0
R1P srcP inP R value={R_s} noisetemp=0 noiseflow=0 dcvar=0 dcvarlot=0
R2N fbN outN R value={R_a} noisetemp=0 noiseflow=0 dcvar={sigma_R^2} dcvarlot={Lot_1}
R2P outP fbP R value={R_a} noisetemp=0 noiseflow=0 dcvar={sigma_R^2} dcvarlot={Lot_1}
R3 fbP fbN R value={R_b} noisetemp=0 noiseflow=0 dcvar={sigma_R^2} dcvarlot=0
R4 outP outN R value={R_L} noisetemp=0 noiseflow=0 dcvar=0 dcvarlot=0
V1N srcN 0 V value=0 noise=0 dc=0 dcvar=0
V1P srcP 0 V value=0 noise=0 dc=0 dcvar=0
X1N inN fbN outN 0 O_dcvar svo={sigma_vo} sio={sigma_io} sib={sigma_ib} iib={I_b}
X1P inP fbP outP 0 O_dcvar svo={sigma_vo} sio={sigma_io} sib={sigma_ib} iib={I_b}
.end